/*
 * punc_interlv_lut - TODO
 *
 * Michael Tetemke Mehari michael.mehari@ugent.be
 */

module punc_interlv_lut
(
  input  wire [3:0] rate,
  input  wire [8:0] idx_i,
  output reg  [8:0] idx_o,
  output reg        punc_o
);

  always @ * begin
    idx_o  = 511;
    punc_o = 1;
	// 6 Mbps
	if(rate == 4'b1011) begin
	  case (idx_i)
		 0: begin idx_o = 0;   punc_o = 0; end
		 1: begin idx_o = 24;  punc_o = 0; end
		 2: begin idx_o = 48;  punc_o = 0; end
		 3: begin idx_o = 72;  punc_o = 0; end
		 4: begin idx_o = 96;  punc_o = 0; end
		 5: begin idx_o = 120; punc_o = 0; end
		 6: begin idx_o = 144; punc_o = 0; end
		 7: begin idx_o = 168; punc_o = 0; end
		 8: begin idx_o = 192; punc_o = 0; end
		 9: begin idx_o = 216; punc_o = 0; end
		10: begin idx_o = 240; punc_o = 0; end
		11: begin idx_o = 264; punc_o = 0; end
		12: begin idx_o = 288; punc_o = 0; end
		13: begin idx_o = 312; punc_o = 0; end
		14: begin idx_o = 336; punc_o = 0; end
		15: begin idx_o = 360; punc_o = 0; end
		16: begin idx_o = 8;   punc_o = 0; end
		17: begin idx_o = 32;  punc_o = 0; end
		18: begin idx_o = 56;  punc_o = 0; end
		19: begin idx_o = 80;  punc_o = 0; end
		20: begin idx_o = 104; punc_o = 0; end
		21: begin idx_o = 128; punc_o = 0; end
		22: begin idx_o = 152; punc_o = 0; end
		23: begin idx_o = 176; punc_o = 0; end
		24: begin idx_o = 200; punc_o = 0; end
		25: begin idx_o = 224; punc_o = 0; end
		26: begin idx_o = 248; punc_o = 0; end
		27: begin idx_o = 272; punc_o = 0; end
		28: begin idx_o = 296; punc_o = 0; end
		29: begin idx_o = 320; punc_o = 0; end
		30: begin idx_o = 344; punc_o = 0; end
		31: begin idx_o = 368; punc_o = 0; end
		32: begin idx_o = 16;  punc_o = 0; end
		33: begin idx_o = 40;  punc_o = 0; end
		34: begin idx_o = 64;  punc_o = 0; end
		35: begin idx_o = 88;  punc_o = 0; end
		36: begin idx_o = 112; punc_o = 0; end
		37: begin idx_o = 136; punc_o = 0; end
		38: begin idx_o = 160; punc_o = 0; end
		39: begin idx_o = 184; punc_o = 0; end
		40: begin idx_o = 208; punc_o = 0; end
		41: begin idx_o = 232; punc_o = 0; end
		42: begin idx_o = 256; punc_o = 0; end
		43: begin idx_o = 280; punc_o = 0; end
		44: begin idx_o = 304; punc_o = 0; end
		45: begin idx_o = 328; punc_o = 0; end
		46: begin idx_o = 352; punc_o = 0; end
		47: begin idx_o = 376; punc_o = 0; end
	  endcase
	end

	// 9 Mbps
	else if(rate == 4'b1111) begin
	  case (idx_i)
		 0: begin idx_o = 0;     punc_o = 0; end
		 1: begin idx_o = 24;    punc_o = 0; end
		 2: begin idx_o = 48;    punc_o = 0; end
		 5: begin idx_o = 72;    punc_o = 0; end
		 6: begin idx_o = 96;    punc_o = 0; end
		 7: begin idx_o = 120;   punc_o = 0; end
		 8: begin idx_o = 144;   punc_o = 0; end
		11: begin idx_o = 168;   punc_o = 0; end
		12: begin idx_o = 192;   punc_o = 0; end
		13: begin idx_o = 216;   punc_o = 0; end
		14: begin idx_o = 240;   punc_o = 0; end
		17: begin idx_o = 264;   punc_o = 0; end
		18: begin idx_o = 288;   punc_o = 0; end
		19: begin idx_o = 312;   punc_o = 0; end
		20: begin idx_o = 336;   punc_o = 0; end
		23: begin idx_o = 360;   punc_o = 0; end
		24: begin idx_o = 8;     punc_o = 0; end
		25: begin idx_o = 32;    punc_o = 0; end
		26: begin idx_o = 56;    punc_o = 0; end
		29: begin idx_o = 80;    punc_o = 0; end
		30: begin idx_o = 104;   punc_o = 0; end
		31: begin idx_o = 128;   punc_o = 0; end
		32: begin idx_o = 152;   punc_o = 0; end
		35: begin idx_o = 176;   punc_o = 0; end
		36: begin idx_o = 200;   punc_o = 0; end
		37: begin idx_o = 224;   punc_o = 0; end
		38: begin idx_o = 248;   punc_o = 0; end
		41: begin idx_o = 272;   punc_o = 0; end
		42: begin idx_o = 296;   punc_o = 0; end
		43: begin idx_o = 320;   punc_o = 0; end
		44: begin idx_o = 344;   punc_o = 0; end
		47: begin idx_o = 368;   punc_o = 0; end
		48: begin idx_o = 16;    punc_o = 0; end
		49: begin idx_o = 40;    punc_o = 0; end
		50: begin idx_o = 64;    punc_o = 0; end
		53: begin idx_o = 88;    punc_o = 0; end
		54: begin idx_o = 112;   punc_o = 0; end
		55: begin idx_o = 136;   punc_o = 0; end
		56: begin idx_o = 160;   punc_o = 0; end
		59: begin idx_o = 184;   punc_o = 0; end
		60: begin idx_o = 208;   punc_o = 0; end
		61: begin idx_o = 232;   punc_o = 0; end
		62: begin idx_o = 256;   punc_o = 0; end
		65: begin idx_o = 280;   punc_o = 0; end
		66: begin idx_o = 304;   punc_o = 0; end
		67: begin idx_o = 328;   punc_o = 0; end
		68: begin idx_o = 352;   punc_o = 0; end
		71: begin idx_o = 376;   punc_o = 0; end
	  endcase
	end

	// 12 Mbps
	else if(rate == 4'b1010) begin
	  case (idx_i)
		 0: begin idx_o = 0;     punc_o = 0; end
		 1: begin idx_o = 24;    punc_o = 0; end
		 2: begin idx_o = 48;    punc_o = 0; end
		 3: begin idx_o = 72;    punc_o = 0; end
		 4: begin idx_o = 96;    punc_o = 0; end
		 5: begin idx_o = 120;   punc_o = 0; end
		 6: begin idx_o = 144;   punc_o = 0; end
		 7: begin idx_o = 168;   punc_o = 0; end
		 8: begin idx_o = 192;   punc_o = 0; end
		 9: begin idx_o = 216;   punc_o = 0; end
		10: begin idx_o = 240;   punc_o = 0; end
		11: begin idx_o = 264;   punc_o = 0; end
		12: begin idx_o = 288;   punc_o = 0; end
		13: begin idx_o = 312;   punc_o = 0; end
		14: begin idx_o = 336;   punc_o = 0; end
		15: begin idx_o = 360;   punc_o = 0; end
		16: begin idx_o = 1;     punc_o = 0; end
		17: begin idx_o = 25;    punc_o = 0; end
		18: begin idx_o = 49;    punc_o = 0; end
		19: begin idx_o = 73;    punc_o = 0; end
		20: begin idx_o = 97;    punc_o = 0; end
		21: begin idx_o = 121;   punc_o = 0; end
		22: begin idx_o = 145;   punc_o = 0; end
		23: begin idx_o = 169;   punc_o = 0; end
		24: begin idx_o = 193;   punc_o = 0; end
		25: begin idx_o = 217;   punc_o = 0; end
		26: begin idx_o = 241;   punc_o = 0; end
		27: begin idx_o = 265;   punc_o = 0; end
		28: begin idx_o = 289;   punc_o = 0; end
		29: begin idx_o = 313;   punc_o = 0; end
		30: begin idx_o = 337;   punc_o = 0; end
		31: begin idx_o = 361;   punc_o = 0; end
		32: begin idx_o = 8;     punc_o = 0; end
		33: begin idx_o = 32;    punc_o = 0; end
		34: begin idx_o = 56;    punc_o = 0; end
		35: begin idx_o = 80;    punc_o = 0; end
		36: begin idx_o = 104;   punc_o = 0; end
		37: begin idx_o = 128;   punc_o = 0; end
		38: begin idx_o = 152;   punc_o = 0; end
		39: begin idx_o = 176;   punc_o = 0; end
		40: begin idx_o = 200;   punc_o = 0; end
		41: begin idx_o = 224;   punc_o = 0; end
		42: begin idx_o = 248;   punc_o = 0; end
		43: begin idx_o = 272;   punc_o = 0; end
		44: begin idx_o = 296;   punc_o = 0; end
		45: begin idx_o = 320;   punc_o = 0; end
		46: begin idx_o = 344;   punc_o = 0; end
		47: begin idx_o = 368;   punc_o = 0; end
		48: begin idx_o = 9;     punc_o = 0; end
		49: begin idx_o = 33;    punc_o = 0; end
		50: begin idx_o = 57;    punc_o = 0; end
		51: begin idx_o = 81;    punc_o = 0; end
		52: begin idx_o = 105;   punc_o = 0; end
		53: begin idx_o = 129;   punc_o = 0; end
		54: begin idx_o = 153;   punc_o = 0; end
		55: begin idx_o = 177;   punc_o = 0; end
		56: begin idx_o = 201;   punc_o = 0; end
		57: begin idx_o = 225;   punc_o = 0; end
		58: begin idx_o = 249;   punc_o = 0; end
		59: begin idx_o = 273;   punc_o = 0; end
		60: begin idx_o = 297;   punc_o = 0; end
		61: begin idx_o = 321;   punc_o = 0; end
		62: begin idx_o = 345;   punc_o = 0; end
		63: begin idx_o = 369;   punc_o = 0; end
		64: begin idx_o = 16;    punc_o = 0; end
		65: begin idx_o = 40;    punc_o = 0; end
		66: begin idx_o = 64;    punc_o = 0; end
		67: begin idx_o = 88;    punc_o = 0; end
		68: begin idx_o = 112;   punc_o = 0; end
		69: begin idx_o = 136;   punc_o = 0; end
		70: begin idx_o = 160;   punc_o = 0; end
		71: begin idx_o = 184;   punc_o = 0; end
		72: begin idx_o = 208;   punc_o = 0; end
		73: begin idx_o = 232;   punc_o = 0; end
		74: begin idx_o = 256;   punc_o = 0; end
		75: begin idx_o = 280;   punc_o = 0; end
		76: begin idx_o = 304;   punc_o = 0; end
		77: begin idx_o = 328;   punc_o = 0; end
		78: begin idx_o = 352;   punc_o = 0; end
		79: begin idx_o = 376;   punc_o = 0; end
		80: begin idx_o = 17;    punc_o = 0; end
		81: begin idx_o = 41;    punc_o = 0; end
		82: begin idx_o = 65;    punc_o = 0; end
		83: begin idx_o = 89;    punc_o = 0; end
		84: begin idx_o = 113;   punc_o = 0; end
		85: begin idx_o = 137;   punc_o = 0; end
		86: begin idx_o = 161;   punc_o = 0; end
		87: begin idx_o = 185;   punc_o = 0; end
		88: begin idx_o = 209;   punc_o = 0; end
		89: begin idx_o = 233;   punc_o = 0; end
		90: begin idx_o = 257;   punc_o = 0; end
		91: begin idx_o = 281;   punc_o = 0; end
		92: begin idx_o = 305;   punc_o = 0; end
		93: begin idx_o = 329;   punc_o = 0; end
		94: begin idx_o = 353;   punc_o = 0; end
		95: begin idx_o = 377;   punc_o = 0; end
	  endcase
	end

	// 18 Mbps
	else if(rate == 4'b1110) begin
	  case (idx_i)
		  0: begin idx_o = 0;     punc_o = 0; end
		  1: begin idx_o = 24;    punc_o = 0; end
		  2: begin idx_o = 48;    punc_o = 0; end
		  5: begin idx_o = 72;    punc_o = 0; end
		  6: begin idx_o = 96;    punc_o = 0; end
		  7: begin idx_o = 120;   punc_o = 0; end
		  8: begin idx_o = 144;   punc_o = 0; end
		 11: begin idx_o = 168;   punc_o = 0; end
		 12: begin idx_o = 192;   punc_o = 0; end
		 13: begin idx_o = 216;   punc_o = 0; end
		 14: begin idx_o = 240;   punc_o = 0; end
		 17: begin idx_o = 264;   punc_o = 0; end
		 18: begin idx_o = 288;   punc_o = 0; end
		 19: begin idx_o = 312;   punc_o = 0; end
		 20: begin idx_o = 336;   punc_o = 0; end
		 23: begin idx_o = 360;   punc_o = 0; end
		 24: begin idx_o = 1;     punc_o = 0; end
		 25: begin idx_o = 25;    punc_o = 0; end
		 26: begin idx_o = 49;    punc_o = 0; end
		 29: begin idx_o = 73;    punc_o = 0; end
		 30: begin idx_o = 97;    punc_o = 0; end
		 31: begin idx_o = 121;   punc_o = 0; end
		 32: begin idx_o = 145;   punc_o = 0; end
		 35: begin idx_o = 169;   punc_o = 0; end
		 36: begin idx_o = 193;   punc_o = 0; end
		 37: begin idx_o = 217;   punc_o = 0; end
		 38: begin idx_o = 241;   punc_o = 0; end
		 41: begin idx_o = 265;   punc_o = 0; end
		 42: begin idx_o = 289;   punc_o = 0; end
		 43: begin idx_o = 313;   punc_o = 0; end
		 44: begin idx_o = 337;   punc_o = 0; end
		 47: begin idx_o = 361;   punc_o = 0; end
		 48: begin idx_o = 8;     punc_o = 0; end
		 49: begin idx_o = 32;    punc_o = 0; end
		 50: begin idx_o = 56;    punc_o = 0; end
		 53: begin idx_o = 80;    punc_o = 0; end
		 54: begin idx_o = 104;   punc_o = 0; end
		 55: begin idx_o = 128;   punc_o = 0; end
		 56: begin idx_o = 152;   punc_o = 0; end
		 59: begin idx_o = 176;   punc_o = 0; end
		 60: begin idx_o = 200;   punc_o = 0; end
		 61: begin idx_o = 224;   punc_o = 0; end
		 62: begin idx_o = 248;   punc_o = 0; end
		 65: begin idx_o = 272;   punc_o = 0; end
		 66: begin idx_o = 296;   punc_o = 0; end
		 67: begin idx_o = 320;   punc_o = 0; end
		 68: begin idx_o = 344;   punc_o = 0; end
		 71: begin idx_o = 368;   punc_o = 0; end
		 72: begin idx_o = 9;     punc_o = 0; end
		 73: begin idx_o = 33;    punc_o = 0; end
		 74: begin idx_o = 57;    punc_o = 0; end
		 77: begin idx_o = 81;    punc_o = 0; end
		 78: begin idx_o = 105;   punc_o = 0; end
		 79: begin idx_o = 129;   punc_o = 0; end
		 80: begin idx_o = 153;   punc_o = 0; end
		 83: begin idx_o = 177;   punc_o = 0; end
		 84: begin idx_o = 201;   punc_o = 0; end
		 85: begin idx_o = 225;   punc_o = 0; end
		 86: begin idx_o = 249;   punc_o = 0; end
		 89: begin idx_o = 273;   punc_o = 0; end
		 90: begin idx_o = 297;   punc_o = 0; end
		 91: begin idx_o = 321;   punc_o = 0; end
		 92: begin idx_o = 345;   punc_o = 0; end
		 95: begin idx_o = 369;   punc_o = 0; end
		 96: begin idx_o = 16;    punc_o = 0; end
		 97: begin idx_o = 40;    punc_o = 0; end
		 98: begin idx_o = 64;    punc_o = 0; end
		101: begin idx_o = 88;    punc_o = 0; end
		102: begin idx_o = 112;   punc_o = 0; end
		103: begin idx_o = 136;   punc_o = 0; end
		104: begin idx_o = 160;   punc_o = 0; end
		107: begin idx_o = 184;   punc_o = 0; end
		108: begin idx_o = 208;   punc_o = 0; end
		109: begin idx_o = 232;   punc_o = 0; end
		110: begin idx_o = 256;   punc_o = 0; end
		113: begin idx_o = 280;   punc_o = 0; end
		114: begin idx_o = 304;   punc_o = 0; end
		115: begin idx_o = 328;   punc_o = 0; end
		116: begin idx_o = 352;   punc_o = 0; end
		119: begin idx_o = 376;   punc_o = 0; end
		120: begin idx_o = 17;    punc_o = 0; end
		121: begin idx_o = 41;    punc_o = 0; end
		122: begin idx_o = 65;    punc_o = 0; end
		125: begin idx_o = 89;    punc_o = 0; end
		126: begin idx_o = 113;   punc_o = 0; end
		127: begin idx_o = 137;   punc_o = 0; end
		128: begin idx_o = 161;   punc_o = 0; end
		131: begin idx_o = 185;   punc_o = 0; end
		132: begin idx_o = 209;   punc_o = 0; end
		133: begin idx_o = 233;   punc_o = 0; end
		134: begin idx_o = 257;   punc_o = 0; end
		137: begin idx_o = 281;   punc_o = 0; end
		138: begin idx_o = 305;   punc_o = 0; end
		139: begin idx_o = 329;   punc_o = 0; end
		140: begin idx_o = 353;   punc_o = 0; end
		143: begin idx_o = 377;   punc_o = 0; end
	  endcase
	end

	// 24 Mbps
	else if(rate == 4'b1001) begin
	  case (idx_i)
		  0: begin idx_o = 0;     punc_o = 0; end
		  1: begin idx_o = 25;    punc_o = 0; end
		  2: begin idx_o = 48;    punc_o = 0; end
		  3: begin idx_o = 73;    punc_o = 0; end
		  4: begin idx_o = 96;    punc_o = 0; end
		  5: begin idx_o = 121;   punc_o = 0; end
		  6: begin idx_o = 144;   punc_o = 0; end
		  7: begin idx_o = 169;   punc_o = 0; end
		  8: begin idx_o = 192;   punc_o = 0; end
		  9: begin idx_o = 217;   punc_o = 0; end
		 10: begin idx_o = 240;   punc_o = 0; end
		 11: begin idx_o = 265;   punc_o = 0; end
		 12: begin idx_o = 288;   punc_o = 0; end
		 13: begin idx_o = 313;   punc_o = 0; end
		 14: begin idx_o = 336;   punc_o = 0; end
		 15: begin idx_o = 361;   punc_o = 0; end
		 16: begin idx_o = 1;     punc_o = 0; end
		 17: begin idx_o = 24;    punc_o = 0; end
		 18: begin idx_o = 49;    punc_o = 0; end
		 19: begin idx_o = 72;    punc_o = 0; end
		 20: begin idx_o = 97;    punc_o = 0; end
		 21: begin idx_o = 120;   punc_o = 0; end
		 22: begin idx_o = 145;   punc_o = 0; end
		 23: begin idx_o = 168;   punc_o = 0; end
		 24: begin idx_o = 193;   punc_o = 0; end
		 25: begin idx_o = 216;   punc_o = 0; end
		 26: begin idx_o = 241;   punc_o = 0; end
		 27: begin idx_o = 264;   punc_o = 0; end
		 28: begin idx_o = 289;   punc_o = 0; end
		 29: begin idx_o = 312;   punc_o = 0; end
		 30: begin idx_o = 337;   punc_o = 0; end
		 31: begin idx_o = 360;   punc_o = 0; end
		 32: begin idx_o = 2;     punc_o = 0; end
		 33: begin idx_o = 27;    punc_o = 0; end
		 34: begin idx_o = 50;    punc_o = 0; end
		 35: begin idx_o = 75;    punc_o = 0; end
		 36: begin idx_o = 98;    punc_o = 0; end
		 37: begin idx_o = 123;   punc_o = 0; end
		 38: begin idx_o = 146;   punc_o = 0; end
		 39: begin idx_o = 171;   punc_o = 0; end
		 40: begin idx_o = 194;   punc_o = 0; end
		 41: begin idx_o = 219;   punc_o = 0; end
		 42: begin idx_o = 242;   punc_o = 0; end
		 43: begin idx_o = 267;   punc_o = 0; end
		 44: begin idx_o = 290;   punc_o = 0; end
		 45: begin idx_o = 315;   punc_o = 0; end
		 46: begin idx_o = 338;   punc_o = 0; end
		 47: begin idx_o = 363;   punc_o = 0; end
		 48: begin idx_o = 3;     punc_o = 0; end
		 49: begin idx_o = 26;    punc_o = 0; end
		 50: begin idx_o = 51;    punc_o = 0; end
		 51: begin idx_o = 74;    punc_o = 0; end
		 52: begin idx_o = 99;    punc_o = 0; end
		 53: begin idx_o = 122;   punc_o = 0; end
		 54: begin idx_o = 147;   punc_o = 0; end
		 55: begin idx_o = 170;   punc_o = 0; end
		 56: begin idx_o = 195;   punc_o = 0; end
		 57: begin idx_o = 218;   punc_o = 0; end
		 58: begin idx_o = 243;   punc_o = 0; end
		 59: begin idx_o = 266;   punc_o = 0; end
		 60: begin idx_o = 291;   punc_o = 0; end
		 61: begin idx_o = 314;   punc_o = 0; end
		 62: begin idx_o = 339;   punc_o = 0; end
		 63: begin idx_o = 362;   punc_o = 0; end
		 64: begin idx_o = 8;     punc_o = 0; end
		 65: begin idx_o = 33;    punc_o = 0; end
		 66: begin idx_o = 56;    punc_o = 0; end
		 67: begin idx_o = 81;    punc_o = 0; end
		 68: begin idx_o = 104;   punc_o = 0; end
		 69: begin idx_o = 129;   punc_o = 0; end
		 70: begin idx_o = 152;   punc_o = 0; end
		 71: begin idx_o = 177;   punc_o = 0; end
		 72: begin idx_o = 200;   punc_o = 0; end
		 73: begin idx_o = 225;   punc_o = 0; end
		 74: begin idx_o = 248;   punc_o = 0; end
		 75: begin idx_o = 273;   punc_o = 0; end
		 76: begin idx_o = 296;   punc_o = 0; end
		 77: begin idx_o = 321;   punc_o = 0; end
		 78: begin idx_o = 344;   punc_o = 0; end
		 79: begin idx_o = 369;   punc_o = 0; end
		 80: begin idx_o = 9;     punc_o = 0; end
		 81: begin idx_o = 32;    punc_o = 0; end
		 82: begin idx_o = 57;    punc_o = 0; end
		 83: begin idx_o = 80;    punc_o = 0; end
		 84: begin idx_o = 105;   punc_o = 0; end
		 85: begin idx_o = 128;   punc_o = 0; end
		 86: begin idx_o = 153;   punc_o = 0; end
		 87: begin idx_o = 176;   punc_o = 0; end
		 88: begin idx_o = 201;   punc_o = 0; end
		 89: begin idx_o = 224;   punc_o = 0; end
		 90: begin idx_o = 249;   punc_o = 0; end
		 91: begin idx_o = 272;   punc_o = 0; end
		 92: begin idx_o = 297;   punc_o = 0; end
		 93: begin idx_o = 320;   punc_o = 0; end
		 94: begin idx_o = 345;   punc_o = 0; end
		 95: begin idx_o = 368;   punc_o = 0; end
		 96: begin idx_o = 10;    punc_o = 0; end
		 97: begin idx_o = 35;    punc_o = 0; end
		 98: begin idx_o = 58;    punc_o = 0; end
		 99: begin idx_o = 83;    punc_o = 0; end
		100: begin idx_o = 106;   punc_o = 0; end
		101: begin idx_o = 131;   punc_o = 0; end
		102: begin idx_o = 154;   punc_o = 0; end
		103: begin idx_o = 179;   punc_o = 0; end
		104: begin idx_o = 202;   punc_o = 0; end
		105: begin idx_o = 227;   punc_o = 0; end
		106: begin idx_o = 250;   punc_o = 0; end
		107: begin idx_o = 275;   punc_o = 0; end
		108: begin idx_o = 298;   punc_o = 0; end
		109: begin idx_o = 323;   punc_o = 0; end
		110: begin idx_o = 346;   punc_o = 0; end
		111: begin idx_o = 371;   punc_o = 0; end
		112: begin idx_o = 11;    punc_o = 0; end
		113: begin idx_o = 34;    punc_o = 0; end
		114: begin idx_o = 59;    punc_o = 0; end
		115: begin idx_o = 82;    punc_o = 0; end
		116: begin idx_o = 107;   punc_o = 0; end
		117: begin idx_o = 130;   punc_o = 0; end
		118: begin idx_o = 155;   punc_o = 0; end
		119: begin idx_o = 178;   punc_o = 0; end
		120: begin idx_o = 203;   punc_o = 0; end
		121: begin idx_o = 226;   punc_o = 0; end
		122: begin idx_o = 251;   punc_o = 0; end
		123: begin idx_o = 274;   punc_o = 0; end
		124: begin idx_o = 299;   punc_o = 0; end
		125: begin idx_o = 322;   punc_o = 0; end
		126: begin idx_o = 347;   punc_o = 0; end
		127: begin idx_o = 370;   punc_o = 0; end
		128: begin idx_o = 16;    punc_o = 0; end
		129: begin idx_o = 41;    punc_o = 0; end
		130: begin idx_o = 64;    punc_o = 0; end
		131: begin idx_o = 89;    punc_o = 0; end
		132: begin idx_o = 112;   punc_o = 0; end
		133: begin idx_o = 137;   punc_o = 0; end
		134: begin idx_o = 160;   punc_o = 0; end
		135: begin idx_o = 185;   punc_o = 0; end
		136: begin idx_o = 208;   punc_o = 0; end
		137: begin idx_o = 233;   punc_o = 0; end
		138: begin idx_o = 256;   punc_o = 0; end
		139: begin idx_o = 281;   punc_o = 0; end
		140: begin idx_o = 304;   punc_o = 0; end
		141: begin idx_o = 329;   punc_o = 0; end
		142: begin idx_o = 352;   punc_o = 0; end
		143: begin idx_o = 377;   punc_o = 0; end
		144: begin idx_o = 17;    punc_o = 0; end
		145: begin idx_o = 40;    punc_o = 0; end
		146: begin idx_o = 65;    punc_o = 0; end
		147: begin idx_o = 88;    punc_o = 0; end
		148: begin idx_o = 113;   punc_o = 0; end
		149: begin idx_o = 136;   punc_o = 0; end
		150: begin idx_o = 161;   punc_o = 0; end
		151: begin idx_o = 184;   punc_o = 0; end
		152: begin idx_o = 209;   punc_o = 0; end
		153: begin idx_o = 232;   punc_o = 0; end
		154: begin idx_o = 257;   punc_o = 0; end
		155: begin idx_o = 280;   punc_o = 0; end
		156: begin idx_o = 305;   punc_o = 0; end
		157: begin idx_o = 328;   punc_o = 0; end
		158: begin idx_o = 353;   punc_o = 0; end
		159: begin idx_o = 376;   punc_o = 0; end
		160: begin idx_o = 18;    punc_o = 0; end
		161: begin idx_o = 43;    punc_o = 0; end
		162: begin idx_o = 66;    punc_o = 0; end
		163: begin idx_o = 91;    punc_o = 0; end
		164: begin idx_o = 114;   punc_o = 0; end
		165: begin idx_o = 139;   punc_o = 0; end
		166: begin idx_o = 162;   punc_o = 0; end
		167: begin idx_o = 187;   punc_o = 0; end
		168: begin idx_o = 210;   punc_o = 0; end
		169: begin idx_o = 235;   punc_o = 0; end
		170: begin idx_o = 258;   punc_o = 0; end
		171: begin idx_o = 283;   punc_o = 0; end
		172: begin idx_o = 306;   punc_o = 0; end
		173: begin idx_o = 331;   punc_o = 0; end
		174: begin idx_o = 354;   punc_o = 0; end
		175: begin idx_o = 379;   punc_o = 0; end
		176: begin idx_o = 19;    punc_o = 0; end
		177: begin idx_o = 42;    punc_o = 0; end
		178: begin idx_o = 67;    punc_o = 0; end
		179: begin idx_o = 90;    punc_o = 0; end
		180: begin idx_o = 115;   punc_o = 0; end
		181: begin idx_o = 138;   punc_o = 0; end
		182: begin idx_o = 163;   punc_o = 0; end
		183: begin idx_o = 186;   punc_o = 0; end
		184: begin idx_o = 211;   punc_o = 0; end
		185: begin idx_o = 234;   punc_o = 0; end
		186: begin idx_o = 259;   punc_o = 0; end
		187: begin idx_o = 282;   punc_o = 0; end
		188: begin idx_o = 307;   punc_o = 0; end
		189: begin idx_o = 330;   punc_o = 0; end
		190: begin idx_o = 355;   punc_o = 0; end
		191: begin idx_o = 378;   punc_o = 0; end
	  endcase
	end

	// 36 Mbps
	else if(rate == 4'b1101) begin
	  case (idx_i)
		  0: begin idx_o = 0;     punc_o = 0; end
		  1: begin idx_o = 25;    punc_o = 0; end
		  2: begin idx_o = 48;    punc_o = 0; end
		  5: begin idx_o = 73;    punc_o = 0; end
		  6: begin idx_o = 96;    punc_o = 0; end
		  7: begin idx_o = 121;   punc_o = 0; end
		  8: begin idx_o = 144;   punc_o = 0; end
		 11: begin idx_o = 169;   punc_o = 0; end
		 12: begin idx_o = 192;   punc_o = 0; end
		 13: begin idx_o = 217;   punc_o = 0; end
		 14: begin idx_o = 240;   punc_o = 0; end
		 17: begin idx_o = 265;   punc_o = 0; end
		 18: begin idx_o = 288;   punc_o = 0; end
		 19: begin idx_o = 313;   punc_o = 0; end
		 20: begin idx_o = 336;   punc_o = 0; end
		 23: begin idx_o = 361;   punc_o = 0; end
		 24: begin idx_o = 1;     punc_o = 0; end
		 25: begin idx_o = 24;    punc_o = 0; end
		 26: begin idx_o = 49;    punc_o = 0; end
		 29: begin idx_o = 72;    punc_o = 0; end
		 30: begin idx_o = 97;    punc_o = 0; end
		 31: begin idx_o = 120;   punc_o = 0; end
		 32: begin idx_o = 145;   punc_o = 0; end
		 35: begin idx_o = 168;   punc_o = 0; end
		 36: begin idx_o = 193;   punc_o = 0; end
		 37: begin idx_o = 216;   punc_o = 0; end
		 38: begin idx_o = 241;   punc_o = 0; end
		 41: begin idx_o = 264;   punc_o = 0; end
		 42: begin idx_o = 289;   punc_o = 0; end
		 43: begin idx_o = 312;   punc_o = 0; end
		 44: begin idx_o = 337;   punc_o = 0; end
		 47: begin idx_o = 360;   punc_o = 0; end
		 48: begin idx_o = 2;     punc_o = 0; end
		 49: begin idx_o = 27;    punc_o = 0; end
		 50: begin idx_o = 50;    punc_o = 0; end
		 53: begin idx_o = 75;    punc_o = 0; end
		 54: begin idx_o = 98;    punc_o = 0; end
		 55: begin idx_o = 123;   punc_o = 0; end
		 56: begin idx_o = 146;   punc_o = 0; end
		 59: begin idx_o = 171;   punc_o = 0; end
		 60: begin idx_o = 194;   punc_o = 0; end
		 61: begin idx_o = 219;   punc_o = 0; end
		 62: begin idx_o = 242;   punc_o = 0; end
		 65: begin idx_o = 267;   punc_o = 0; end
		 66: begin idx_o = 290;   punc_o = 0; end
		 67: begin idx_o = 315;   punc_o = 0; end
		 68: begin idx_o = 338;   punc_o = 0; end
		 71: begin idx_o = 363;   punc_o = 0; end
		 72: begin idx_o = 3;     punc_o = 0; end
		 73: begin idx_o = 26;    punc_o = 0; end
		 74: begin idx_o = 51;    punc_o = 0; end
		 77: begin idx_o = 74;    punc_o = 0; end
		 78: begin idx_o = 99;    punc_o = 0; end
		 79: begin idx_o = 122;   punc_o = 0; end
		 80: begin idx_o = 147;   punc_o = 0; end
		 83: begin idx_o = 170;   punc_o = 0; end
		 84: begin idx_o = 195;   punc_o = 0; end
		 85: begin idx_o = 218;   punc_o = 0; end
		 86: begin idx_o = 243;   punc_o = 0; end
		 89: begin idx_o = 266;   punc_o = 0; end
		 90: begin idx_o = 291;   punc_o = 0; end
		 91: begin idx_o = 314;   punc_o = 0; end
		 92: begin idx_o = 339;   punc_o = 0; end
		 95: begin idx_o = 362;   punc_o = 0; end
		 96: begin idx_o = 8;     punc_o = 0; end
		 97: begin idx_o = 33;    punc_o = 0; end
		 98: begin idx_o = 56;    punc_o = 0; end
		101: begin idx_o = 81;    punc_o = 0; end
		102: begin idx_o = 104;   punc_o = 0; end
		103: begin idx_o = 129;   punc_o = 0; end
		104: begin idx_o = 152;   punc_o = 0; end
		107: begin idx_o = 177;   punc_o = 0; end
		108: begin idx_o = 200;   punc_o = 0; end
		109: begin idx_o = 225;   punc_o = 0; end
		110: begin idx_o = 248;   punc_o = 0; end
		113: begin idx_o = 273;   punc_o = 0; end
		114: begin idx_o = 296;   punc_o = 0; end
		115: begin idx_o = 321;   punc_o = 0; end
		116: begin idx_o = 344;   punc_o = 0; end
		119: begin idx_o = 369;   punc_o = 0; end
		120: begin idx_o = 9;     punc_o = 0; end
		121: begin idx_o = 32;    punc_o = 0; end
		122: begin idx_o = 57;    punc_o = 0; end
		125: begin idx_o = 80;    punc_o = 0; end
		126: begin idx_o = 105;   punc_o = 0; end
		127: begin idx_o = 128;   punc_o = 0; end
		128: begin idx_o = 153;   punc_o = 0; end
		131: begin idx_o = 176;   punc_o = 0; end
		132: begin idx_o = 201;   punc_o = 0; end
		133: begin idx_o = 224;   punc_o = 0; end
		134: begin idx_o = 249;   punc_o = 0; end
		137: begin idx_o = 272;   punc_o = 0; end
		138: begin idx_o = 297;   punc_o = 0; end
		139: begin idx_o = 320;   punc_o = 0; end
		140: begin idx_o = 345;   punc_o = 0; end
		143: begin idx_o = 368;   punc_o = 0; end
		144: begin idx_o = 10;    punc_o = 0; end
		145: begin idx_o = 35;    punc_o = 0; end
		146: begin idx_o = 58;    punc_o = 0; end
		149: begin idx_o = 83;    punc_o = 0; end
		150: begin idx_o = 106;   punc_o = 0; end
		151: begin idx_o = 131;   punc_o = 0; end
		152: begin idx_o = 154;   punc_o = 0; end
		155: begin idx_o = 179;   punc_o = 0; end
		156: begin idx_o = 202;   punc_o = 0; end
		157: begin idx_o = 227;   punc_o = 0; end
		158: begin idx_o = 250;   punc_o = 0; end
		161: begin idx_o = 275;   punc_o = 0; end
		162: begin idx_o = 298;   punc_o = 0; end
		163: begin idx_o = 323;   punc_o = 0; end
		164: begin idx_o = 346;   punc_o = 0; end
		167: begin idx_o = 371;   punc_o = 0; end
		168: begin idx_o = 11;    punc_o = 0; end
		169: begin idx_o = 34;    punc_o = 0; end
		170: begin idx_o = 59;    punc_o = 0; end
		173: begin idx_o = 82;    punc_o = 0; end
		174: begin idx_o = 107;   punc_o = 0; end
		175: begin idx_o = 130;   punc_o = 0; end
		176: begin idx_o = 155;   punc_o = 0; end
		179: begin idx_o = 178;   punc_o = 0; end
		180: begin idx_o = 203;   punc_o = 0; end
		181: begin idx_o = 226;   punc_o = 0; end
		182: begin idx_o = 251;   punc_o = 0; end
		185: begin idx_o = 274;   punc_o = 0; end
		186: begin idx_o = 299;   punc_o = 0; end
		187: begin idx_o = 322;   punc_o = 0; end
		188: begin idx_o = 347;   punc_o = 0; end
		191: begin idx_o = 370;   punc_o = 0; end
		192: begin idx_o = 16;    punc_o = 0; end
		193: begin idx_o = 41;    punc_o = 0; end
		194: begin idx_o = 64;    punc_o = 0; end
		197: begin idx_o = 89;    punc_o = 0; end
		198: begin idx_o = 112;   punc_o = 0; end
		199: begin idx_o = 137;   punc_o = 0; end
		200: begin idx_o = 160;   punc_o = 0; end
		203: begin idx_o = 185;   punc_o = 0; end
		204: begin idx_o = 208;   punc_o = 0; end
		205: begin idx_o = 233;   punc_o = 0; end
		206: begin idx_o = 256;   punc_o = 0; end
		209: begin idx_o = 281;   punc_o = 0; end
		210: begin idx_o = 304;   punc_o = 0; end
		211: begin idx_o = 329;   punc_o = 0; end
		212: begin idx_o = 352;   punc_o = 0; end
		215: begin idx_o = 377;   punc_o = 0; end
		216: begin idx_o = 17;    punc_o = 0; end
		217: begin idx_o = 40;    punc_o = 0; end
		218: begin idx_o = 65;    punc_o = 0; end
		221: begin idx_o = 88;    punc_o = 0; end
		222: begin idx_o = 113;   punc_o = 0; end
		223: begin idx_o = 136;   punc_o = 0; end
		224: begin idx_o = 161;   punc_o = 0; end
		227: begin idx_o = 184;   punc_o = 0; end
		228: begin idx_o = 209;   punc_o = 0; end
		229: begin idx_o = 232;   punc_o = 0; end
		230: begin idx_o = 257;   punc_o = 0; end
		233: begin idx_o = 280;   punc_o = 0; end
		234: begin idx_o = 305;   punc_o = 0; end
		235: begin idx_o = 328;   punc_o = 0; end
		236: begin idx_o = 353;   punc_o = 0; end
		239: begin idx_o = 376;   punc_o = 0; end
		240: begin idx_o = 18;    punc_o = 0; end
		241: begin idx_o = 43;    punc_o = 0; end
		242: begin idx_o = 66;    punc_o = 0; end
		245: begin idx_o = 91;    punc_o = 0; end
		246: begin idx_o = 114;   punc_o = 0; end
		247: begin idx_o = 139;   punc_o = 0; end
		248: begin idx_o = 162;   punc_o = 0; end
		251: begin idx_o = 187;   punc_o = 0; end
		252: begin idx_o = 210;   punc_o = 0; end
		253: begin idx_o = 235;   punc_o = 0; end
		254: begin idx_o = 258;   punc_o = 0; end
		257: begin idx_o = 283;   punc_o = 0; end
		258: begin idx_o = 306;   punc_o = 0; end
		259: begin idx_o = 331;   punc_o = 0; end
		260: begin idx_o = 354;   punc_o = 0; end
		263: begin idx_o = 379;   punc_o = 0; end
		264: begin idx_o = 19;    punc_o = 0; end
		265: begin idx_o = 42;    punc_o = 0; end
		266: begin idx_o = 67;    punc_o = 0; end
		269: begin idx_o = 90;    punc_o = 0; end
		270: begin idx_o = 115;   punc_o = 0; end
		271: begin idx_o = 138;   punc_o = 0; end
		272: begin idx_o = 163;   punc_o = 0; end
		275: begin idx_o = 186;   punc_o = 0; end
		276: begin idx_o = 211;   punc_o = 0; end
		277: begin idx_o = 234;   punc_o = 0; end
		278: begin idx_o = 259;   punc_o = 0; end
		281: begin idx_o = 282;   punc_o = 0; end
		282: begin idx_o = 307;   punc_o = 0; end
		283: begin idx_o = 330;   punc_o = 0; end
		284: begin idx_o = 355;   punc_o = 0; end
		287: begin idx_o = 378;   punc_o = 0; end        
	  endcase
	end

	// 48 Mbps
	else if(rate == 4'b1000) begin
	  case (idx_i)
		  0: begin idx_o = 0;     punc_o = 0; end
		  1: begin idx_o = 26;    punc_o = 0; end
		  2: begin idx_o = 49;    punc_o = 0; end
		  4: begin idx_o = 72;    punc_o = 0; end
		  5: begin idx_o = 98;    punc_o = 0; end
		  6: begin idx_o = 121;   punc_o = 0; end
		  8: begin idx_o = 144;   punc_o = 0; end
		  9: begin idx_o = 170;   punc_o = 0; end
		 10: begin idx_o = 193;   punc_o = 0; end
		 12: begin idx_o = 216;   punc_o = 0; end
		 13: begin idx_o = 242;   punc_o = 0; end
		 14: begin idx_o = 265;   punc_o = 0; end
		 16: begin idx_o = 288;   punc_o = 0; end
		 17: begin idx_o = 314;   punc_o = 0; end
		 18: begin idx_o = 337;   punc_o = 0; end
		 20: begin idx_o = 360;   punc_o = 0; end
		 21: begin idx_o = 1;     punc_o = 0; end
		 22: begin idx_o = 24;    punc_o = 0; end
		 24: begin idx_o = 50;    punc_o = 0; end
		 25: begin idx_o = 73;    punc_o = 0; end
		 26: begin idx_o = 96;    punc_o = 0; end
		 28: begin idx_o = 122;   punc_o = 0; end
		 29: begin idx_o = 145;   punc_o = 0; end
		 30: begin idx_o = 168;   punc_o = 0; end
		 32: begin idx_o = 194;   punc_o = 0; end
		 33: begin idx_o = 217;   punc_o = 0; end
		 34: begin idx_o = 240;   punc_o = 0; end
		 36: begin idx_o = 266;   punc_o = 0; end
		 37: begin idx_o = 289;   punc_o = 0; end
		 38: begin idx_o = 312;   punc_o = 0; end
		 40: begin idx_o = 338;   punc_o = 0; end
		 41: begin idx_o = 361;   punc_o = 0; end
		 42: begin idx_o = 2;     punc_o = 0; end
		 44: begin idx_o = 25;    punc_o = 0; end
		 45: begin idx_o = 48;    punc_o = 0; end
		 46: begin idx_o = 74;    punc_o = 0; end
		 48: begin idx_o = 97;    punc_o = 0; end
		 49: begin idx_o = 120;   punc_o = 0; end
		 50: begin idx_o = 146;   punc_o = 0; end
		 52: begin idx_o = 169;   punc_o = 0; end
		 53: begin idx_o = 192;   punc_o = 0; end
		 54: begin idx_o = 218;   punc_o = 0; end
		 56: begin idx_o = 241;   punc_o = 0; end
		 57: begin idx_o = 264;   punc_o = 0; end
		 58: begin idx_o = 290;   punc_o = 0; end
		 60: begin idx_o = 313;   punc_o = 0; end
		 61: begin idx_o = 336;   punc_o = 0; end
		 62: begin idx_o = 362;   punc_o = 0; end
		 64: begin idx_o = 3;     punc_o = 0; end
		 65: begin idx_o = 29;    punc_o = 0; end
		 66: begin idx_o = 52;    punc_o = 0; end
		 68: begin idx_o = 75;    punc_o = 0; end
		 69: begin idx_o = 101;   punc_o = 0; end
		 70: begin idx_o = 124;   punc_o = 0; end
		 72: begin idx_o = 147;   punc_o = 0; end
		 73: begin idx_o = 173;   punc_o = 0; end
		 74: begin idx_o = 196;   punc_o = 0; end
		 76: begin idx_o = 219;   punc_o = 0; end
		 77: begin idx_o = 245;   punc_o = 0; end
		 78: begin idx_o = 268;   punc_o = 0; end
		 80: begin idx_o = 291;   punc_o = 0; end
		 81: begin idx_o = 317;   punc_o = 0; end
		 82: begin idx_o = 340;   punc_o = 0; end
		 84: begin idx_o = 363;   punc_o = 0; end
		 85: begin idx_o = 4;     punc_o = 0; end
		 86: begin idx_o = 27;    punc_o = 0; end
		 88: begin idx_o = 53;    punc_o = 0; end
		 89: begin idx_o = 76;    punc_o = 0; end
		 90: begin idx_o = 99;    punc_o = 0; end
		 92: begin idx_o = 125;   punc_o = 0; end
		 93: begin idx_o = 148;   punc_o = 0; end
		 94: begin idx_o = 171;   punc_o = 0; end
		 96: begin idx_o = 197;   punc_o = 0; end
		 97: begin idx_o = 220;   punc_o = 0; end
		 98: begin idx_o = 243;   punc_o = 0; end
		100: begin idx_o = 269;   punc_o = 0; end
		101: begin idx_o = 292;   punc_o = 0; end
		102: begin idx_o = 315;   punc_o = 0; end
		104: begin idx_o = 341;   punc_o = 0; end
		105: begin idx_o = 364;   punc_o = 0; end
		106: begin idx_o = 5;     punc_o = 0; end
		108: begin idx_o = 28;    punc_o = 0; end
		109: begin idx_o = 51;    punc_o = 0; end
		110: begin idx_o = 77;    punc_o = 0; end
		112: begin idx_o = 100;   punc_o = 0; end
		113: begin idx_o = 123;   punc_o = 0; end
		114: begin idx_o = 149;   punc_o = 0; end
		116: begin idx_o = 172;   punc_o = 0; end
		117: begin idx_o = 195;   punc_o = 0; end
		118: begin idx_o = 221;   punc_o = 0; end
		120: begin idx_o = 244;   punc_o = 0; end
		121: begin idx_o = 267;   punc_o = 0; end
		122: begin idx_o = 293;   punc_o = 0; end
		124: begin idx_o = 316;   punc_o = 0; end
		125: begin idx_o = 339;   punc_o = 0; end
		126: begin idx_o = 365;   punc_o = 0; end
		128: begin idx_o = 8;     punc_o = 0; end
		129: begin idx_o = 34;    punc_o = 0; end
		130: begin idx_o = 57;    punc_o = 0; end
		132: begin idx_o = 80;    punc_o = 0; end
		133: begin idx_o = 106;   punc_o = 0; end
		134: begin idx_o = 129;   punc_o = 0; end
		136: begin idx_o = 152;   punc_o = 0; end
		137: begin idx_o = 178;   punc_o = 0; end
		138: begin idx_o = 201;   punc_o = 0; end
		140: begin idx_o = 224;   punc_o = 0; end
		141: begin idx_o = 250;   punc_o = 0; end
		142: begin idx_o = 273;   punc_o = 0; end
		144: begin idx_o = 296;   punc_o = 0; end
		145: begin idx_o = 322;   punc_o = 0; end
		146: begin idx_o = 345;   punc_o = 0; end
		148: begin idx_o = 368;   punc_o = 0; end
		149: begin idx_o = 9;     punc_o = 0; end
		150: begin idx_o = 32;    punc_o = 0; end
		152: begin idx_o = 58;    punc_o = 0; end
		153: begin idx_o = 81;    punc_o = 0; end
		154: begin idx_o = 104;   punc_o = 0; end
		156: begin idx_o = 130;   punc_o = 0; end
		157: begin idx_o = 153;   punc_o = 0; end
		158: begin idx_o = 176;   punc_o = 0; end
		160: begin idx_o = 202;   punc_o = 0; end
		161: begin idx_o = 225;   punc_o = 0; end
		162: begin idx_o = 248;   punc_o = 0; end
		164: begin idx_o = 274;   punc_o = 0; end
		165: begin idx_o = 297;   punc_o = 0; end
		166: begin idx_o = 320;   punc_o = 0; end
		168: begin idx_o = 346;   punc_o = 0; end
		169: begin idx_o = 369;   punc_o = 0; end
		170: begin idx_o = 10;    punc_o = 0; end
		172: begin idx_o = 33;    punc_o = 0; end
		173: begin idx_o = 56;    punc_o = 0; end
		174: begin idx_o = 82;    punc_o = 0; end
		176: begin idx_o = 105;   punc_o = 0; end
		177: begin idx_o = 128;   punc_o = 0; end
		178: begin idx_o = 154;   punc_o = 0; end
		180: begin idx_o = 177;   punc_o = 0; end
		181: begin idx_o = 200;   punc_o = 0; end
		182: begin idx_o = 226;   punc_o = 0; end
		184: begin idx_o = 249;   punc_o = 0; end
		185: begin idx_o = 272;   punc_o = 0; end
		186: begin idx_o = 298;   punc_o = 0; end
		188: begin idx_o = 321;   punc_o = 0; end
		189: begin idx_o = 344;   punc_o = 0; end
		190: begin idx_o = 370;   punc_o = 0; end
		192: begin idx_o = 11;    punc_o = 0; end
		193: begin idx_o = 37;    punc_o = 0; end
		194: begin idx_o = 60;    punc_o = 0; end
		196: begin idx_o = 83;    punc_o = 0; end
		197: begin idx_o = 109;   punc_o = 0; end
		198: begin idx_o = 132;   punc_o = 0; end
		200: begin idx_o = 155;   punc_o = 0; end
		201: begin idx_o = 181;   punc_o = 0; end
		202: begin idx_o = 204;   punc_o = 0; end
		204: begin idx_o = 227;   punc_o = 0; end
		205: begin idx_o = 253;   punc_o = 0; end
		206: begin idx_o = 276;   punc_o = 0; end
		208: begin idx_o = 299;   punc_o = 0; end
		209: begin idx_o = 325;   punc_o = 0; end
		210: begin idx_o = 348;   punc_o = 0; end
		212: begin idx_o = 371;   punc_o = 0; end
		213: begin idx_o = 12;    punc_o = 0; end
		214: begin idx_o = 35;    punc_o = 0; end
		216: begin idx_o = 61;    punc_o = 0; end
		217: begin idx_o = 84;    punc_o = 0; end
		218: begin idx_o = 107;   punc_o = 0; end
		220: begin idx_o = 133;   punc_o = 0; end
		221: begin idx_o = 156;   punc_o = 0; end
		222: begin idx_o = 179;   punc_o = 0; end
		224: begin idx_o = 205;   punc_o = 0; end
		225: begin idx_o = 228;   punc_o = 0; end
		226: begin idx_o = 251;   punc_o = 0; end
		228: begin idx_o = 277;   punc_o = 0; end
		229: begin idx_o = 300;   punc_o = 0; end
		230: begin idx_o = 323;   punc_o = 0; end
		232: begin idx_o = 349;   punc_o = 0; end
		233: begin idx_o = 372;   punc_o = 0; end
		234: begin idx_o = 13;    punc_o = 0; end
		236: begin idx_o = 36;    punc_o = 0; end
		237: begin idx_o = 59;    punc_o = 0; end
		238: begin idx_o = 85;    punc_o = 0; end
		240: begin idx_o = 108;   punc_o = 0; end
		241: begin idx_o = 131;   punc_o = 0; end
		242: begin idx_o = 157;   punc_o = 0; end
		244: begin idx_o = 180;   punc_o = 0; end
		245: begin idx_o = 203;   punc_o = 0; end
		246: begin idx_o = 229;   punc_o = 0; end
		248: begin idx_o = 252;   punc_o = 0; end
		249: begin idx_o = 275;   punc_o = 0; end
		250: begin idx_o = 301;   punc_o = 0; end
		252: begin idx_o = 324;   punc_o = 0; end
		253: begin idx_o = 347;   punc_o = 0; end
		254: begin idx_o = 373;   punc_o = 0; end
		256: begin idx_o = 16;    punc_o = 0; end
		257: begin idx_o = 42;    punc_o = 0; end
		258: begin idx_o = 65;    punc_o = 0; end
		260: begin idx_o = 88;    punc_o = 0; end
		261: begin idx_o = 114;   punc_o = 0; end
		262: begin idx_o = 137;   punc_o = 0; end
		264: begin idx_o = 160;   punc_o = 0; end
		265: begin idx_o = 186;   punc_o = 0; end
		266: begin idx_o = 209;   punc_o = 0; end
		268: begin idx_o = 232;   punc_o = 0; end
		269: begin idx_o = 258;   punc_o = 0; end
		270: begin idx_o = 281;   punc_o = 0; end
		272: begin idx_o = 304;   punc_o = 0; end
		273: begin idx_o = 330;   punc_o = 0; end
		274: begin idx_o = 353;   punc_o = 0; end
		276: begin idx_o = 376;   punc_o = 0; end
		277: begin idx_o = 17;    punc_o = 0; end
		278: begin idx_o = 40;    punc_o = 0; end
		280: begin idx_o = 66;    punc_o = 0; end
		281: begin idx_o = 89;    punc_o = 0; end
		282: begin idx_o = 112;   punc_o = 0; end
		284: begin idx_o = 138;   punc_o = 0; end
		285: begin idx_o = 161;   punc_o = 0; end
		286: begin idx_o = 184;   punc_o = 0; end
		288: begin idx_o = 210;   punc_o = 0; end
		289: begin idx_o = 233;   punc_o = 0; end
		290: begin idx_o = 256;   punc_o = 0; end
		292: begin idx_o = 282;   punc_o = 0; end
		293: begin idx_o = 305;   punc_o = 0; end
		294: begin idx_o = 328;   punc_o = 0; end
		296: begin idx_o = 354;   punc_o = 0; end
		297: begin idx_o = 377;   punc_o = 0; end
		298: begin idx_o = 18;    punc_o = 0; end
		300: begin idx_o = 41;    punc_o = 0; end
		301: begin idx_o = 64;    punc_o = 0; end
		302: begin idx_o = 90;    punc_o = 0; end
		304: begin idx_o = 113;   punc_o = 0; end
		305: begin idx_o = 136;   punc_o = 0; end
		306: begin idx_o = 162;   punc_o = 0; end
		308: begin idx_o = 185;   punc_o = 0; end
		309: begin idx_o = 208;   punc_o = 0; end
		310: begin idx_o = 234;   punc_o = 0; end
		312: begin idx_o = 257;   punc_o = 0; end
		313: begin idx_o = 280;   punc_o = 0; end
		314: begin idx_o = 306;   punc_o = 0; end
		316: begin idx_o = 329;   punc_o = 0; end
		317: begin idx_o = 352;   punc_o = 0; end
		318: begin idx_o = 378;   punc_o = 0; end
		320: begin idx_o = 19;    punc_o = 0; end
		321: begin idx_o = 45;    punc_o = 0; end
		322: begin idx_o = 68;    punc_o = 0; end
		324: begin idx_o = 91;    punc_o = 0; end
		325: begin idx_o = 117;   punc_o = 0; end
		326: begin idx_o = 140;   punc_o = 0; end
		328: begin idx_o = 163;   punc_o = 0; end
		329: begin idx_o = 189;   punc_o = 0; end
		330: begin idx_o = 212;   punc_o = 0; end
		332: begin idx_o = 235;   punc_o = 0; end
		333: begin idx_o = 261;   punc_o = 0; end
		334: begin idx_o = 284;   punc_o = 0; end
		336: begin idx_o = 307;   punc_o = 0; end
		337: begin idx_o = 333;   punc_o = 0; end
		338: begin idx_o = 356;   punc_o = 0; end
		340: begin idx_o = 379;   punc_o = 0; end
		341: begin idx_o = 20;    punc_o = 0; end
		342: begin idx_o = 43;    punc_o = 0; end
		344: begin idx_o = 69;    punc_o = 0; end
		345: begin idx_o = 92;    punc_o = 0; end
		346: begin idx_o = 115;   punc_o = 0; end
		348: begin idx_o = 141;   punc_o = 0; end
		349: begin idx_o = 164;   punc_o = 0; end
		350: begin idx_o = 187;   punc_o = 0; end
		352: begin idx_o = 213;   punc_o = 0; end
		353: begin idx_o = 236;   punc_o = 0; end
		354: begin idx_o = 259;   punc_o = 0; end
		356: begin idx_o = 285;   punc_o = 0; end
		357: begin idx_o = 308;   punc_o = 0; end
		358: begin idx_o = 331;   punc_o = 0; end
		360: begin idx_o = 357;   punc_o = 0; end
		361: begin idx_o = 380;   punc_o = 0; end
		362: begin idx_o = 21;    punc_o = 0; end
		364: begin idx_o = 44;    punc_o = 0; end
		365: begin idx_o = 67;    punc_o = 0; end
		366: begin idx_o = 93;    punc_o = 0; end
		368: begin idx_o = 116;   punc_o = 0; end
		369: begin idx_o = 139;   punc_o = 0; end
		370: begin idx_o = 165;   punc_o = 0; end
		372: begin idx_o = 188;   punc_o = 0; end
		373: begin idx_o = 211;   punc_o = 0; end
		374: begin idx_o = 237;   punc_o = 0; end
		376: begin idx_o = 260;   punc_o = 0; end
		377: begin idx_o = 283;   punc_o = 0; end
		378: begin idx_o = 309;   punc_o = 0; end
		380: begin idx_o = 332;   punc_o = 0; end
		381: begin idx_o = 355;   punc_o = 0; end
		382: begin idx_o = 381;   punc_o = 0; end
	  endcase
	end

	// 54 Mbps
	else if(rate == 4'b1100) begin
	  case (idx_i)
          0: begin idx_o = 0;     punc_o = 0; end
		  1: begin idx_o = 26;    punc_o = 0; end
		  2: begin idx_o = 49;    punc_o = 0; end
		  5: begin idx_o = 72;    punc_o = 0; end
		  6: begin idx_o = 98;    punc_o = 0; end
		  7: begin idx_o = 121;   punc_o = 0; end
		  8: begin idx_o = 144;   punc_o = 0; end
		 11: begin idx_o = 170;   punc_o = 0; end
		 12: begin idx_o = 193;   punc_o = 0; end
		 13: begin idx_o = 216;   punc_o = 0; end
		 14: begin idx_o = 242;   punc_o = 0; end
		 17: begin idx_o = 265;   punc_o = 0; end
		 18: begin idx_o = 288;   punc_o = 0; end
		 19: begin idx_o = 314;   punc_o = 0; end
		 20: begin idx_o = 337;   punc_o = 0; end
		 23: begin idx_o = 360;   punc_o = 0; end
		 24: begin idx_o = 1;     punc_o = 0; end
		 25: begin idx_o = 24;    punc_o = 0; end
		 26: begin idx_o = 50;    punc_o = 0; end
		 29: begin idx_o = 73;    punc_o = 0; end
		 30: begin idx_o = 96;    punc_o = 0; end
		 31: begin idx_o = 122;   punc_o = 0; end
		 32: begin idx_o = 145;   punc_o = 0; end
		 35: begin idx_o = 168;   punc_o = 0; end
		 36: begin idx_o = 194;   punc_o = 0; end
		 37: begin idx_o = 217;   punc_o = 0; end
		 38: begin idx_o = 240;   punc_o = 0; end
		 41: begin idx_o = 266;   punc_o = 0; end
		 42: begin idx_o = 289;   punc_o = 0; end
		 43: begin idx_o = 312;   punc_o = 0; end
		 44: begin idx_o = 338;   punc_o = 0; end
		 47: begin idx_o = 361;   punc_o = 0; end
		 48: begin idx_o = 2;     punc_o = 0; end
		 49: begin idx_o = 25;    punc_o = 0; end
		 50: begin idx_o = 48;    punc_o = 0; end
		 53: begin idx_o = 74;    punc_o = 0; end
		 54: begin idx_o = 97;    punc_o = 0; end
		 55: begin idx_o = 120;   punc_o = 0; end
		 56: begin idx_o = 146;   punc_o = 0; end
		 59: begin idx_o = 169;   punc_o = 0; end
		 60: begin idx_o = 192;   punc_o = 0; end
		 61: begin idx_o = 218;   punc_o = 0; end
		 62: begin idx_o = 241;   punc_o = 0; end
		 65: begin idx_o = 264;   punc_o = 0; end
		 66: begin idx_o = 290;   punc_o = 0; end
		 67: begin idx_o = 313;   punc_o = 0; end
		 68: begin idx_o = 336;   punc_o = 0; end
		 71: begin idx_o = 362;   punc_o = 0; end
		 72: begin idx_o = 3;     punc_o = 0; end
		 73: begin idx_o = 29;    punc_o = 0; end
		 74: begin idx_o = 52;    punc_o = 0; end
		 77: begin idx_o = 75;    punc_o = 0; end
		 78: begin idx_o = 101;   punc_o = 0; end
		 79: begin idx_o = 124;   punc_o = 0; end
		 80: begin idx_o = 147;   punc_o = 0; end
		 83: begin idx_o = 173;   punc_o = 0; end
		 84: begin idx_o = 196;   punc_o = 0; end
		 85: begin idx_o = 219;   punc_o = 0; end
		 86: begin idx_o = 245;   punc_o = 0; end
		 89: begin idx_o = 268;   punc_o = 0; end
		 90: begin idx_o = 291;   punc_o = 0; end
		 91: begin idx_o = 317;   punc_o = 0; end
		 92: begin idx_o = 340;   punc_o = 0; end
		 95: begin idx_o = 363;   punc_o = 0; end
		 96: begin idx_o = 4;     punc_o = 0; end
		 97: begin idx_o = 27;    punc_o = 0; end
		 98: begin idx_o = 53;    punc_o = 0; end
		101: begin idx_o = 76;    punc_o = 0; end
		102: begin idx_o = 99;    punc_o = 0; end
		103: begin idx_o = 125;   punc_o = 0; end
		104: begin idx_o = 148;   punc_o = 0; end
		107: begin idx_o = 171;   punc_o = 0; end
		108: begin idx_o = 197;   punc_o = 0; end
		109: begin idx_o = 220;   punc_o = 0; end
		110: begin idx_o = 243;   punc_o = 0; end
		113: begin idx_o = 269;   punc_o = 0; end
		114: begin idx_o = 292;   punc_o = 0; end
		115: begin idx_o = 315;   punc_o = 0; end
		116: begin idx_o = 341;   punc_o = 0; end
		119: begin idx_o = 364;   punc_o = 0; end
		120: begin idx_o = 5;     punc_o = 0; end
		121: begin idx_o = 28;    punc_o = 0; end
		122: begin idx_o = 51;    punc_o = 0; end
		125: begin idx_o = 77;    punc_o = 0; end
		126: begin idx_o = 100;   punc_o = 0; end
		127: begin idx_o = 123;   punc_o = 0; end
		128: begin idx_o = 149;   punc_o = 0; end
		131: begin idx_o = 172;   punc_o = 0; end
		132: begin idx_o = 195;   punc_o = 0; end
		133: begin idx_o = 221;   punc_o = 0; end
		134: begin idx_o = 244;   punc_o = 0; end
		137: begin idx_o = 267;   punc_o = 0; end
		138: begin idx_o = 293;   punc_o = 0; end
		139: begin idx_o = 316;   punc_o = 0; end
		140: begin idx_o = 339;   punc_o = 0; end
		143: begin idx_o = 365;   punc_o = 0; end
		144: begin idx_o = 8;     punc_o = 0; end
		145: begin idx_o = 34;    punc_o = 0; end
		146: begin idx_o = 57;    punc_o = 0; end
		149: begin idx_o = 80;    punc_o = 0; end
		150: begin idx_o = 106;   punc_o = 0; end
		151: begin idx_o = 129;   punc_o = 0; end
		152: begin idx_o = 152;   punc_o = 0; end
		155: begin idx_o = 178;   punc_o = 0; end
		156: begin idx_o = 201;   punc_o = 0; end
		157: begin idx_o = 224;   punc_o = 0; end
		158: begin idx_o = 250;   punc_o = 0; end
		161: begin idx_o = 273;   punc_o = 0; end
		162: begin idx_o = 296;   punc_o = 0; end
		163: begin idx_o = 322;   punc_o = 0; end
		164: begin idx_o = 345;   punc_o = 0; end
		167: begin idx_o = 368;   punc_o = 0; end
		168: begin idx_o = 9;     punc_o = 0; end
		169: begin idx_o = 32;    punc_o = 0; end
		170: begin idx_o = 58;    punc_o = 0; end
		173: begin idx_o = 81;    punc_o = 0; end
		174: begin idx_o = 104;   punc_o = 0; end
		175: begin idx_o = 130;   punc_o = 0; end
		176: begin idx_o = 153;   punc_o = 0; end
		179: begin idx_o = 176;   punc_o = 0; end
		180: begin idx_o = 202;   punc_o = 0; end
		181: begin idx_o = 225;   punc_o = 0; end
		182: begin idx_o = 248;   punc_o = 0; end
		185: begin idx_o = 274;   punc_o = 0; end
		186: begin idx_o = 297;   punc_o = 0; end
		187: begin idx_o = 320;   punc_o = 0; end
		188: begin idx_o = 346;   punc_o = 0; end
		191: begin idx_o = 369;   punc_o = 0; end
		192: begin idx_o = 10;    punc_o = 0; end
		193: begin idx_o = 33;    punc_o = 0; end
		194: begin idx_o = 56;    punc_o = 0; end
		197: begin idx_o = 82;    punc_o = 0; end
		198: begin idx_o = 105;   punc_o = 0; end
		199: begin idx_o = 128;   punc_o = 0; end
		200: begin idx_o = 154;   punc_o = 0; end
		203: begin idx_o = 177;   punc_o = 0; end
		204: begin idx_o = 200;   punc_o = 0; end
		205: begin idx_o = 226;   punc_o = 0; end
		206: begin idx_o = 249;   punc_o = 0; end
		209: begin idx_o = 272;   punc_o = 0; end
		210: begin idx_o = 298;   punc_o = 0; end
		211: begin idx_o = 321;   punc_o = 0; end
		212: begin idx_o = 344;   punc_o = 0; end
		215: begin idx_o = 370;   punc_o = 0; end
		216: begin idx_o = 11;    punc_o = 0; end
		217: begin idx_o = 37;    punc_o = 0; end
		218: begin idx_o = 60;    punc_o = 0; end
		221: begin idx_o = 83;    punc_o = 0; end
		222: begin idx_o = 109;   punc_o = 0; end
		223: begin idx_o = 132;   punc_o = 0; end
		224: begin idx_o = 155;   punc_o = 0; end
		227: begin idx_o = 181;   punc_o = 0; end
		228: begin idx_o = 204;   punc_o = 0; end
		229: begin idx_o = 227;   punc_o = 0; end
		230: begin idx_o = 253;   punc_o = 0; end
		233: begin idx_o = 276;   punc_o = 0; end
		234: begin idx_o = 299;   punc_o = 0; end
		235: begin idx_o = 325;   punc_o = 0; end
		236: begin idx_o = 348;   punc_o = 0; end
		239: begin idx_o = 371;   punc_o = 0; end
		240: begin idx_o = 12;    punc_o = 0; end
		241: begin idx_o = 35;    punc_o = 0; end
		242: begin idx_o = 61;    punc_o = 0; end
		245: begin idx_o = 84;    punc_o = 0; end
		246: begin idx_o = 107;   punc_o = 0; end
		247: begin idx_o = 133;   punc_o = 0; end
		248: begin idx_o = 156;   punc_o = 0; end
		251: begin idx_o = 179;   punc_o = 0; end
		252: begin idx_o = 205;   punc_o = 0; end
		253: begin idx_o = 228;   punc_o = 0; end
		254: begin idx_o = 251;   punc_o = 0; end
		257: begin idx_o = 277;   punc_o = 0; end
		258: begin idx_o = 300;   punc_o = 0; end
		259: begin idx_o = 323;   punc_o = 0; end
		260: begin idx_o = 349;   punc_o = 0; end
		263: begin idx_o = 372;   punc_o = 0; end
		264: begin idx_o = 13;    punc_o = 0; end
		265: begin idx_o = 36;    punc_o = 0; end
		266: begin idx_o = 59;    punc_o = 0; end
		269: begin idx_o = 85;    punc_o = 0; end
		270: begin idx_o = 108;   punc_o = 0; end
		271: begin idx_o = 131;   punc_o = 0; end
		272: begin idx_o = 157;   punc_o = 0; end
		275: begin idx_o = 180;   punc_o = 0; end
		276: begin idx_o = 203;   punc_o = 0; end
		277: begin idx_o = 229;   punc_o = 0; end
		278: begin idx_o = 252;   punc_o = 0; end
		281: begin idx_o = 275;   punc_o = 0; end
		282: begin idx_o = 301;   punc_o = 0; end
		283: begin idx_o = 324;   punc_o = 0; end
		284: begin idx_o = 347;   punc_o = 0; end
		287: begin idx_o = 373;   punc_o = 0; end
		288: begin idx_o = 16;    punc_o = 0; end
		289: begin idx_o = 42;    punc_o = 0; end
		290: begin idx_o = 65;    punc_o = 0; end
		293: begin idx_o = 88;    punc_o = 0; end
		294: begin idx_o = 114;   punc_o = 0; end
		295: begin idx_o = 137;   punc_o = 0; end
		296: begin idx_o = 160;   punc_o = 0; end
		299: begin idx_o = 186;   punc_o = 0; end
		300: begin idx_o = 209;   punc_o = 0; end
		301: begin idx_o = 232;   punc_o = 0; end
		302: begin idx_o = 258;   punc_o = 0; end
		305: begin idx_o = 281;   punc_o = 0; end
		306: begin idx_o = 304;   punc_o = 0; end
		307: begin idx_o = 330;   punc_o = 0; end
		308: begin idx_o = 353;   punc_o = 0; end
		311: begin idx_o = 376;   punc_o = 0; end
		312: begin idx_o = 17;    punc_o = 0; end
		313: begin idx_o = 40;    punc_o = 0; end
		314: begin idx_o = 66;    punc_o = 0; end
		317: begin idx_o = 89;    punc_o = 0; end
		318: begin idx_o = 112;   punc_o = 0; end
		319: begin idx_o = 138;   punc_o = 0; end
		320: begin idx_o = 161;   punc_o = 0; end
		323: begin idx_o = 184;   punc_o = 0; end
		324: begin idx_o = 210;   punc_o = 0; end
		325: begin idx_o = 233;   punc_o = 0; end
		326: begin idx_o = 256;   punc_o = 0; end
		329: begin idx_o = 282;   punc_o = 0; end
		330: begin idx_o = 305;   punc_o = 0; end
		331: begin idx_o = 328;   punc_o = 0; end
		332: begin idx_o = 354;   punc_o = 0; end
		335: begin idx_o = 377;   punc_o = 0; end
		336: begin idx_o = 18;    punc_o = 0; end
		337: begin idx_o = 41;    punc_o = 0; end
		338: begin idx_o = 64;    punc_o = 0; end
		341: begin idx_o = 90;    punc_o = 0; end
		342: begin idx_o = 113;   punc_o = 0; end
		343: begin idx_o = 136;   punc_o = 0; end
		344: begin idx_o = 162;   punc_o = 0; end
		347: begin idx_o = 185;   punc_o = 0; end
		348: begin idx_o = 208;   punc_o = 0; end
		349: begin idx_o = 234;   punc_o = 0; end
		350: begin idx_o = 257;   punc_o = 0; end
		353: begin idx_o = 280;   punc_o = 0; end
		354: begin idx_o = 306;   punc_o = 0; end
		355: begin idx_o = 329;   punc_o = 0; end
		356: begin idx_o = 352;   punc_o = 0; end
		359: begin idx_o = 378;   punc_o = 0; end
		360: begin idx_o = 19;    punc_o = 0; end
		361: begin idx_o = 45;    punc_o = 0; end
		362: begin idx_o = 68;    punc_o = 0; end
		365: begin idx_o = 91;    punc_o = 0; end
		366: begin idx_o = 117;   punc_o = 0; end
		367: begin idx_o = 140;   punc_o = 0; end
		368: begin idx_o = 163;   punc_o = 0; end
		371: begin idx_o = 189;   punc_o = 0; end
		372: begin idx_o = 212;   punc_o = 0; end
		373: begin idx_o = 235;   punc_o = 0; end
		374: begin idx_o = 261;   punc_o = 0; end
		377: begin idx_o = 284;   punc_o = 0; end
		378: begin idx_o = 307;   punc_o = 0; end
		379: begin idx_o = 333;   punc_o = 0; end
		380: begin idx_o = 356;   punc_o = 0; end
		383: begin idx_o = 379;   punc_o = 0; end
		384: begin idx_o = 20;    punc_o = 0; end
		385: begin idx_o = 43;    punc_o = 0; end
		386: begin idx_o = 69;    punc_o = 0; end
		389: begin idx_o = 92;    punc_o = 0; end
		390: begin idx_o = 115;   punc_o = 0; end
		391: begin idx_o = 141;   punc_o = 0; end
		392: begin idx_o = 164;   punc_o = 0; end
		395: begin idx_o = 187;   punc_o = 0; end
		396: begin idx_o = 213;   punc_o = 0; end
		397: begin idx_o = 236;   punc_o = 0; end
		398: begin idx_o = 259;   punc_o = 0; end
		401: begin idx_o = 285;   punc_o = 0; end
		402: begin idx_o = 308;   punc_o = 0; end
		403: begin idx_o = 331;   punc_o = 0; end
		404: begin idx_o = 357;   punc_o = 0; end
		407: begin idx_o = 380;   punc_o = 0; end
		408: begin idx_o = 21;    punc_o = 0; end
		409: begin idx_o = 44;    punc_o = 0; end
		410: begin idx_o = 67;    punc_o = 0; end
		413: begin idx_o = 93;    punc_o = 0; end
		414: begin idx_o = 116;   punc_o = 0; end
		415: begin idx_o = 139;   punc_o = 0; end
		416: begin idx_o = 165;   punc_o = 0; end
		419: begin idx_o = 188;   punc_o = 0; end
		420: begin idx_o = 211;   punc_o = 0; end
		421: begin idx_o = 237;   punc_o = 0; end
		422: begin idx_o = 260;   punc_o = 0; end
		425: begin idx_o = 283;   punc_o = 0; end
		426: begin idx_o = 309;   punc_o = 0; end
		427: begin idx_o = 332;   punc_o = 0; end
		428: begin idx_o = 355;   punc_o = 0; end
		431: begin idx_o = 381;   punc_o = 0; end
	  endcase
	end
end
endmodule
